//
// tinybootrom:  bootrom to load applications over i2c
//    for source, see hexloader.as
//
// convert from binary using something like
//    xxd -c2 -a  hexloader.bin |\
//        awk '{printf "         10'\''h%03x: dataout_d = 16'\''h%s;\n", 0x180+NR-1,$2}'

// using global clock and output enable uses no extra resources
// over a combinatorial ROM
//
module tinybootrom(address,dataout);
   input[9:0]   address;
   output[15:0]   dataout;

   // following the idiom in the xilinx guide
   reg  [15:0]  dataout_d;

   assign dataout  = dataout_d ;

   always @ (*)
     begin
       case ( address )
         10'h180: dataout_d = 16'h00a2; // ldx#
         10'h181: dataout_d = 16'h0004;
         10'h182: dataout_d = 16'h009b; // txd special!
         10'h183: dataout_d = 16'h00a2; // ldx#
         10'h184: dataout_d = 16'h0011; //      17
         10'h185: dataout_d = 16'h00a9; // lda#
         10'h186: dataout_d = 16'hf10f; //
         10'h187: dataout_d = 16'h002a; // rol a
         10'h188: dataout_d = 16'h00ca; // dex
         10'h189: dataout_d = 16'h00d0; // bne
         10'h18a: dataout_d = 16'hfffc; //     fc
         10'h18b: dataout_d = 16'h00a2; // ldx#
         10'h18c: dataout_d = 16'h0011; //
         10'h18d: dataout_d = 16'h006a; // ror a
         10'h18e: dataout_d = 16'h00ca; // dex
         10'h18f: dataout_d = 16'h00d0; // bne
         10'h190: dataout_d = 16'hfffc; //     fc
         10'h191: dataout_d = 16'h00a2; // ldx#
         10'h192: dataout_d = 16'h0011; //
         10'h193: dataout_d = 16'h000a; // asl a
         10'h194: dataout_d = 16'h00ca; // dex
         10'h195: dataout_d = 16'h00d0; // bne
         10'h196: dataout_d = 16'hfffc; //     fc
         10'h197: dataout_d = 16'h00a2; // ldx#
         10'h198: dataout_d = 16'h0011; //
         10'h199: dataout_d = 16'h00a9; // lda#
         10'h19a: dataout_d = 16'hF105; //
         10'h19b: dataout_d = 16'h004a; // lsr a
         10'h19c: dataout_d = 16'h00ca; // dex
         10'h19d: dataout_d = 16'h00d0; // bne
         10'h19e: dataout_d = 16'hfffc; //     fc
         10'h19f: dataout_d = 16'h00a2; // ldx#
         10'h1a0: dataout_d = 16'h0011; //
         10'h1a1: dataout_d = 16'h00a9; // lda#
         10'h1a2: dataout_d = 16'h71F5; //
         10'h1a3: dataout_d = 16'h004a; // lsr a
         10'h1a4: dataout_d = 16'h00ca; // dex
         10'h1a5: dataout_d = 16'h00d0; // bne
         10'h1a6: dataout_d = 16'hfffc; //     fc
         10'h1a7: dataout_d = 16'h00f0; // beq
         10'h1a8: dataout_d = 16'hfffe; //     fe (here)
         10'h1a9: dataout_d = 16'h00ea; // nop
         10'h1aa: dataout_d = 16'h00ea; // nop
         10'h1ab: dataout_d = 16'h00ea; // nop
         10'h1ac: dataout_d = 16'h00ea; // nop
         10'h1ad: dataout_d = 16'h00f0; // beq
         10'h1ae: dataout_d = 16'hfffe; //     fe (here)
         10'h1af: dataout_d = 16'h00ea; // nop
         10'h1b0: dataout_d = 16'h006f;
         10'h1b1: dataout_d = 16'h0064;
         10'h1b2: dataout_d = 16'h0065;
         10'h1b3: dataout_d = 16'h0020;
         10'h1b4: dataout_d = 16'h0069;
         10'h1b5: dataout_d = 16'h006a;
         10'h1b6: dataout_d = 16'h0020;
         10'h1b7: dataout_d = 16'h0076;
         10'h1b8: dataout_d = 16'h0061;
         10'h1b9: dataout_d = 16'h0072;
         10'h1ba: dataout_d = 16'h0069;
         10'h1bb: dataout_d = 16'h0061;
         10'h1bc: dataout_d = 16'h006a;
         10'h1bd: dataout_d = 16'h0074;
         10'h1be: dataout_d = 16'h0020;
         10'h1bf: dataout_d = 16'h0049;
         10'h1c0: dataout_d = 16'h006a;
         10'h1c1: dataout_d = 16'h0074;
         10'h1c2: dataout_d = 16'h0065;
         10'h1c3: dataout_d = 16'h006c;
         10'h1c4: dataout_d = 16'h0020;
         10'h1c5: dataout_d = 16'h0048;
         10'h1c6: dataout_d = 16'h0065;
         10'h1c7: dataout_d = 16'h0078;
         10'h1c8: dataout_d = 16'h0020;
         10'h1c9: dataout_d = 16'h0066;
         10'h1ca: dataout_d = 16'h006f;
         10'h1cb: dataout_d = 16'h0072;
         10'h1cc: dataout_d = 16'h006d;
         10'h1cd: dataout_d = 16'h0061;
         10'h1ce: dataout_d = 16'h0074;
         10'h1cf: dataout_d = 16'h0020;
         10'h1d0: dataout_d = 16'h0061;
         10'h1d1: dataout_d = 16'h0074;
         10'h1d2: dataout_d = 16'h0020;
         10'h1d3: dataout_d = 16'h0031;
         10'h1d4: dataout_d = 16'h0039;
         10'h1d5: dataout_d = 16'h0032;
         10'h1d6: dataout_d = 16'h0030;
         10'h1d7: dataout_d = 16'h0030;
         10'h1d8: dataout_d = 16'h002c;
         10'h1d9: dataout_d = 16'h006a;
         10'h1da: dataout_d = 16'h002c;
         10'h1db: dataout_d = 16'h0038;
         10'h1dc: dataout_d = 16'h002c;
         10'h1dd: dataout_d = 16'h0031;
         10'h1de: dataout_d = 16'h0020;
         10'h1df: dataout_d = 16'h002d;
         10'h1e0: dataout_d = 16'h003a;
         10'h1e1: dataout_d = 16'h000d;
         10'h1e2: dataout_d = 16'h000a;
         10'h1e3: dataout_d = 16'h0000;
         10'h1e4: dataout_d = 16'h0020;
         10'h1e5: dataout_d = 16'hff35;
         10'h1e6: dataout_d = 16'hffff;
         10'h1e7: dataout_d = 16'h00c9;
         10'h1e8: dataout_d = 16'h003b;
         10'h1e9: dataout_d = 16'h00d0;
         10'h1ea: dataout_d = 16'hfff9;
         10'h1eb: dataout_d = 16'h00a9;
         10'h1ec: dataout_d = 16'h0000;
         10'h1ed: dataout_d = 16'h0085;
         10'h1ee: dataout_d = 16'h008b;
         10'h1ef: dataout_d = 16'h0020;
         10'h1f0: dataout_d = 16'hff08;
         10'h1f1: dataout_d = 16'hffff;
         10'h1f2: dataout_d = 16'h0085;
         10'h1f3: dataout_d = 16'h0087;
         10'h1f4: dataout_d = 16'h0020;
         10'h1f5: dataout_d = 16'hfef5;
         10'h1f6: dataout_d = 16'hffff;
         10'h1f7: dataout_d = 16'h0085;
         10'h1f8: dataout_d = 16'h0088;
         10'h1f9: dataout_d = 16'h0020;
         10'h1fa: dataout_d = 16'hff08;
         10'h1fb: dataout_d = 16'hffff;
         10'h1fc: dataout_d = 16'h0085;
         10'h1fd: dataout_d = 16'h008a;
         10'h1fe: dataout_d = 16'h00d0;
         10'h1ff: dataout_d = 16'h0027;
         10'h200: dataout_d = 16'h00a6;
         10'h201: dataout_d = 16'h0087;
         10'h202: dataout_d = 16'h00a0;
         10'h203: dataout_d = 16'h0000;
         10'h204: dataout_d = 16'h0020;
         10'h205: dataout_d = 16'hfef5;
         10'h206: dataout_d = 16'hffff;
         10'h207: dataout_d = 16'h0091;
         10'h208: dataout_d = 16'h0088;
         10'h209: dataout_d = 16'h00c8;
         10'h20a: dataout_d = 16'h00ca;
         10'h20b: dataout_d = 16'h00ca;
         10'h20c: dataout_d = 16'h00d0;
         10'h20d: dataout_d = 16'hfff6;
         10'h20e: dataout_d = 16'h0020;
         10'h20f: dataout_d = 16'hff08;
         10'h210: dataout_d = 16'hffff;
         10'h211: dataout_d = 16'h00a5;
         10'h212: dataout_d = 16'h008b;
         10'h213: dataout_d = 16'h00d0;
         10'h214: dataout_d = 16'h0008;
         10'h215: dataout_d = 16'h00a9;
         10'h216: dataout_d = 16'h0023;
         10'h217: dataout_d = 16'h008d;
         10'h218: dataout_d = 16'hfff9;
         10'h219: dataout_d = 16'hfffa;
         10'h21a: dataout_d = 16'h004c;
         10'h21b: dataout_d = 16'hfde4;
         10'h21c: dataout_d = 16'hffff;
         10'h21d: dataout_d = 16'h00a9;
         10'h21e: dataout_d = 16'h0046;
         10'h21f: dataout_d = 16'h0085;
         10'h220: dataout_d = 16'h008c;
         10'h221: dataout_d = 16'h0020;
         10'h222: dataout_d = 16'hff97;
         10'h223: dataout_d = 16'hffff;
         10'h224: dataout_d = 16'h004c;
         10'h225: dataout_d = 16'hfde4;
         10'h226: dataout_d = 16'hffff;
         10'h227: dataout_d = 16'h00c9;
         10'h228: dataout_d = 16'h0001;
         10'h229: dataout_d = 16'h00f0;
         10'h22a: dataout_d = 16'h0031;
         10'h22b: dataout_d = 16'h0020;
         10'h22c: dataout_d = 16'hff5d;
         10'h22d: dataout_d = 16'hffff;
         10'h22e: dataout_d = 16'h000d;
         10'h22f: dataout_d = 16'h000a;
         10'h230: dataout_d = 16'h000d;
         10'h231: dataout_d = 16'h000a;
         10'h232: dataout_d = 16'h0055;
         10'h233: dataout_d = 16'h006a;
         10'h234: dataout_d = 16'h006b;
         10'h235: dataout_d = 16'h006a;
         10'h236: dataout_d = 16'h006f;
         10'h237: dataout_d = 16'h0077;
         10'h238: dataout_d = 16'h006a;
         10'h239: dataout_d = 16'h0020;
         10'h23a: dataout_d = 16'h0072;
         10'h23b: dataout_d = 16'h0065;
         10'h23c: dataout_d = 16'h0063;
         10'h23d: dataout_d = 16'h006f;
         10'h23e: dataout_d = 16'h0072;
         10'h23f: dataout_d = 16'h0064;
         10'h240: dataout_d = 16'h0020;
         10'h241: dataout_d = 16'h0074;
         10'h242: dataout_d = 16'h0079;
         10'h243: dataout_d = 16'h0070;
         10'h244: dataout_d = 16'h0065;
         10'h245: dataout_d = 16'h0020;
         10'h246: dataout_d = 16'h0024;
         10'h247: dataout_d = 16'h0000;
         10'h248: dataout_d = 16'h00a5;
         10'h249: dataout_d = 16'h008a;
         10'h24a: dataout_d = 16'h0085;
         10'h24b: dataout_d = 16'h008c;
         10'h24c: dataout_d = 16'h0020;
         10'h24d: dataout_d = 16'hff84;
         10'h24e: dataout_d = 16'hffff;
         10'h24f: dataout_d = 16'h00a9;
         10'h250: dataout_d = 16'h000d;
         10'h251: dataout_d = 16'h0020;
         10'h252: dataout_d = 16'hff97;
         10'h253: dataout_d = 16'hffff;
         10'h254: dataout_d = 16'h00a9;
         10'h255: dataout_d = 16'h000a;
         10'h256: dataout_d = 16'h0020;
         10'h257: dataout_d = 16'hff97;
         10'h258: dataout_d = 16'hffff;
         10'h259: dataout_d = 16'h004c;
         10'h25a: dataout_d = 16'hfde4;
         10'h25b: dataout_d = 16'hffff;
         10'h25c: dataout_d = 16'h0020;
         10'h25d: dataout_d = 16'hff08;
         10'h25e: dataout_d = 16'hffff;
         10'h25f: dataout_d = 16'h00a5;
         10'h260: dataout_d = 16'h008b;
         10'h261: dataout_d = 16'h00f0;
         10'h262: dataout_d = 16'h0021;
         10'h263: dataout_d = 16'h0020;
         10'h264: dataout_d = 16'hff5d;
         10'h265: dataout_d = 16'hffff;
         10'h266: dataout_d = 16'h000d;
         10'h267: dataout_d = 16'h000a;
         10'h268: dataout_d = 16'h000d;
         10'h269: dataout_d = 16'h000a;
         10'h26a: dataout_d = 16'h0042;
         10'h26b: dataout_d = 16'h0061;
         10'h26c: dataout_d = 16'h0064;
         10'h26d: dataout_d = 16'h0020;
         10'h26e: dataout_d = 16'h0072;
         10'h26f: dataout_d = 16'h0065;
         10'h270: dataout_d = 16'h0063;
         10'h271: dataout_d = 16'h006f;
         10'h272: dataout_d = 16'h0072;
         10'h273: dataout_d = 16'h0064;
         10'h274: dataout_d = 16'h0020;
         10'h275: dataout_d = 16'h0063;
         10'h276: dataout_d = 16'h0068;
         10'h277: dataout_d = 16'h0065;
         10'h278: dataout_d = 16'h0063;
         10'h279: dataout_d = 16'h006b;
         10'h27a: dataout_d = 16'h0073;
         10'h27b: dataout_d = 16'h0075;
         10'h27c: dataout_d = 16'h006d;
         10'h27d: dataout_d = 16'h0021;
         10'h27e: dataout_d = 16'h000d;
         10'h27f: dataout_d = 16'h000a;
         10'h280: dataout_d = 16'h0000;
         10'h281: dataout_d = 16'h004c;
         10'h282: dataout_d = 16'hfd95;
         10'h283: dataout_d = 16'hffff;
         10'h284: dataout_d = 16'h00a5;
         10'h285: dataout_d = 16'h008c;
         10'h286: dataout_d = 16'h00f0;
         10'h287: dataout_d = 16'h0027;
         10'h288: dataout_d = 16'h0020;
         10'h289: dataout_d = 16'hff5d;
         10'h28a: dataout_d = 16'hffff;
         10'h28b: dataout_d = 16'h000d;
         10'h28c: dataout_d = 16'h000a;
         10'h28d: dataout_d = 16'h000d;
         10'h28e: dataout_d = 16'h000a;
         10'h28f: dataout_d = 16'h0044;
         10'h290: dataout_d = 16'h006f;
         10'h291: dataout_d = 16'h0077;
         10'h292: dataout_d = 16'h006a;
         10'h293: dataout_d = 16'h006c;
         10'h294: dataout_d = 16'h006f;
         10'h295: dataout_d = 16'h0061;
         10'h296: dataout_d = 16'h0064;
         10'h297: dataout_d = 16'h0020;
         10'h298: dataout_d = 16'h0046;
         10'h299: dataout_d = 16'h0061;
         10'h29a: dataout_d = 16'h0069;
         10'h29b: dataout_d = 16'h006c;
         10'h29c: dataout_d = 16'h0065;
         10'h29d: dataout_d = 16'h0064;
         10'h29e: dataout_d = 16'h000d;
         10'h29f: dataout_d = 16'h000a;
         10'h2a0: dataout_d = 16'h0041;
         10'h2a1: dataout_d = 16'h0062;
         10'h2a2: dataout_d = 16'h006f;
         10'h2a3: dataout_d = 16'h0072;
         10'h2a4: dataout_d = 16'h0074;
         10'h2a5: dataout_d = 16'h0069;
         10'h2a6: dataout_d = 16'h006a;
         10'h2a7: dataout_d = 16'h0067;
         10'h2a8: dataout_d = 16'h0021;
         10'h2a9: dataout_d = 16'h000d;
         10'h2aa: dataout_d = 16'h000a;
         10'h2ab: dataout_d = 16'h0000;
         10'h2ac: dataout_d = 16'h004c;
         10'h2ad: dataout_d = 16'hfd95;
         10'h2ae: dataout_d = 16'hffff;
         10'h2af: dataout_d = 16'h0020;
         10'h2b0: dataout_d = 16'hff5d;
         10'h2b1: dataout_d = 16'hffff;
         10'h2b2: dataout_d = 16'h000d;
         10'h2b3: dataout_d = 16'h000a;
         10'h2b4: dataout_d = 16'h000d;
         10'h2b5: dataout_d = 16'h000a;
         10'h2b6: dataout_d = 16'h0044;
         10'h2b7: dataout_d = 16'h006f;
         10'h2b8: dataout_d = 16'h0077;
         10'h2b9: dataout_d = 16'h006a;
         10'h2ba: dataout_d = 16'h006c;
         10'h2bb: dataout_d = 16'h006f;
         10'h2bc: dataout_d = 16'h0061;
         10'h2bd: dataout_d = 16'h0064;
         10'h2be: dataout_d = 16'h0020;
         10'h2bf: dataout_d = 16'h0053;
         10'h2c0: dataout_d = 16'h0075;
         10'h2c1: dataout_d = 16'h0063;
         10'h2c2: dataout_d = 16'h0063;
         10'h2c3: dataout_d = 16'h0065;
         10'h2c4: dataout_d = 16'h0073;
         10'h2c5: dataout_d = 16'h0073;
         10'h2c6: dataout_d = 16'h0066;
         10'h2c7: dataout_d = 16'h0075;
         10'h2c8: dataout_d = 16'h006c;
         10'h2c9: dataout_d = 16'h0021;
         10'h2ca: dataout_d = 16'h000d;
         10'h2cb: dataout_d = 16'h000a;
         10'h2cc: dataout_d = 16'h004a;
         10'h2cd: dataout_d = 16'h0075;
         10'h2ce: dataout_d = 16'h006d;
         10'h2cf: dataout_d = 16'h0070;
         10'h2d0: dataout_d = 16'h0069;
         10'h2d1: dataout_d = 16'h006a;
         10'h2d2: dataout_d = 16'h0067;
         10'h2d3: dataout_d = 16'h0020;
         10'h2d4: dataout_d = 16'h0074;
         10'h2d5: dataout_d = 16'h006f;
         10'h2d6: dataout_d = 16'h0020;
         10'h2d7: dataout_d = 16'h006c;
         10'h2d8: dataout_d = 16'h006f;
         10'h2d9: dataout_d = 16'h0063;
         10'h2da: dataout_d = 16'h0061;
         10'h2db: dataout_d = 16'h0074;
         10'h2dc: dataout_d = 16'h0069;
         10'h2dd: dataout_d = 16'h006f;
         10'h2de: dataout_d = 16'h006a;
         10'h2df: dataout_d = 16'h0020;
         10'h2e0: dataout_d = 16'h0024;
         10'h2e1: dataout_d = 16'h0000;
         10'h2e2: dataout_d = 16'h00a9;
         10'h2e3: dataout_d = 16'h0002;
         10'h2e4: dataout_d = 16'h0020;
         10'h2e5: dataout_d = 16'hff84;
         10'h2e6: dataout_d = 16'hffff;
         10'h2e7: dataout_d = 16'h00a9;
         10'h2e8: dataout_d = 16'h0000;
         10'h2e9: dataout_d = 16'h0020;
         10'h2ea: dataout_d = 16'hff84;
         10'h2eb: dataout_d = 16'hffff;
         10'h2ec: dataout_d = 16'h0020;
         10'h2ed: dataout_d = 16'hff5d;
         10'h2ee: dataout_d = 16'hffff;
         10'h2ef: dataout_d = 16'h000d;
         10'h2f0: dataout_d = 16'h000a;
         10'h2f1: dataout_d = 16'h0000;
         10'h2f2: dataout_d = 16'h004c;
         10'h2f3: dataout_d = 16'h0200;
         10'h2f4: dataout_d = 16'h0000;
         10'h2f5: dataout_d = 16'h0020;
         10'h2f6: dataout_d = 16'hff08;
         10'h2f7: dataout_d = 16'hffff;
         10'h2f8: dataout_d = 16'h000a;
         10'h2f9: dataout_d = 16'h000a;
         10'h2fa: dataout_d = 16'h000a;
         10'h2fb: dataout_d = 16'h000a;
         10'h2fc: dataout_d = 16'h000a;
         10'h2fd: dataout_d = 16'h000a;
         10'h2fe: dataout_d = 16'h000a;
         10'h2ff: dataout_d = 16'h000a;
         10'h300: dataout_d = 16'h0085;
         10'h301: dataout_d = 16'h008a;
         10'h302: dataout_d = 16'h0020;
         10'h303: dataout_d = 16'hff08;
         10'h304: dataout_d = 16'hffff;
         10'h305: dataout_d = 16'h0005;
         10'h306: dataout_d = 16'h008a;
         10'h307: dataout_d = 16'h0060;
         10'h308: dataout_d = 16'h0020;
         10'h309: dataout_d = 16'hff35;
         10'h30a: dataout_d = 16'hffff;
         10'h30b: dataout_d = 16'h0020;
         10'h30c: dataout_d = 16'hff2a;
         10'h30d: dataout_d = 16'hffff;
         10'h30e: dataout_d = 16'h000a;
         10'h30f: dataout_d = 16'h000a;
         10'h310: dataout_d = 16'h000a;
         10'h311: dataout_d = 16'h000a;
         10'h312: dataout_d = 16'h0029;
         10'h313: dataout_d = 16'h00f0;
         10'h314: dataout_d = 16'h0085;
         10'h315: dataout_d = 16'h008d;
         10'h316: dataout_d = 16'h0020;
         10'h317: dataout_d = 16'hff35;
         10'h318: dataout_d = 16'hffff;
         10'h319: dataout_d = 16'h0020;
         10'h31a: dataout_d = 16'hff2a;
         10'h31b: dataout_d = 16'hffff;
         10'h31c: dataout_d = 16'h0005;
         10'h31d: dataout_d = 16'h008d;
         10'h31e: dataout_d = 16'h0085;
         10'h31f: dataout_d = 16'h008d;
         10'h320: dataout_d = 16'h0018;
         10'h321: dataout_d = 16'h0065;
         10'h322: dataout_d = 16'h008b;
         10'h323: dataout_d = 16'h0029;
         10'h324: dataout_d = 16'h00ff;
         10'h325: dataout_d = 16'h0085;
         10'h326: dataout_d = 16'h008b;
         10'h327: dataout_d = 16'h00a5;
         10'h328: dataout_d = 16'h008d;
         10'h329: dataout_d = 16'h0060;
         10'h32a: dataout_d = 16'h00c9;
         10'h32b: dataout_d = 16'h003a;
         10'h32c: dataout_d = 16'h0090;
         10'h32d: dataout_d = 16'h0002;
         10'h32e: dataout_d = 16'h00e9;
         10'h32f: dataout_d = 16'h0008;
         10'h330: dataout_d = 16'h00e9;
         10'h331: dataout_d = 16'h002f;
         10'h332: dataout_d = 16'h0029;
         10'h333: dataout_d = 16'h000f;
         10'h334: dataout_d = 16'h0060;
         10'h335: dataout_d = 16'h008a;
         10'h336: dataout_d = 16'h0048;
         10'h337: dataout_d = 16'h00ad;
         10'h338: dataout_d = 16'hfff8;
         10'h339: dataout_d = 16'hfffa;
         10'h33a: dataout_d = 16'h004a;
         10'h33b: dataout_d = 16'h00b0;
         10'h33c: dataout_d = 16'h0017;
         10'h33d: dataout_d = 16'h004a;
         10'h33e: dataout_d = 16'h0090;
         10'h33f: dataout_d = 16'hfff7;
         10'h340: dataout_d = 16'h00a6;
         10'h341: dataout_d = 16'h0082;
         10'h342: dataout_d = 16'h00e4;
         10'h343: dataout_d = 16'h0081;
         10'h344: dataout_d = 16'h00f0;
         10'h345: dataout_d = 16'hfff1;
         10'h346: dataout_d = 16'h00b5;
         10'h347: dataout_d = 16'h0041;
         10'h348: dataout_d = 16'h008d;
         10'h349: dataout_d = 16'hfff9;
         10'h34a: dataout_d = 16'hfffa;
         10'h34b: dataout_d = 16'h00e8;
         10'h34c: dataout_d = 16'h008a;
         10'h34d: dataout_d = 16'h0029;
         10'h34e: dataout_d = 16'h003f;
         10'h34f: dataout_d = 16'h0085;
         10'h350: dataout_d = 16'h0082;
         10'h351: dataout_d = 16'h004c;
         10'h352: dataout_d = 16'hff37;
         10'h353: dataout_d = 16'hffff;
         10'h354: dataout_d = 16'h0068;
         10'h355: dataout_d = 16'h00aa;
         10'h356: dataout_d = 16'h00ad;
         10'h357: dataout_d = 16'hfff9;
         10'h358: dataout_d = 16'hfffa;
         10'h359: dataout_d = 16'h008d;
         10'h35a: dataout_d = 16'h0000;
         10'h35b: dataout_d = 16'hfffd;
         10'h35c: dataout_d = 16'h0060;
         10'h35d: dataout_d = 16'h0084;
         10'h35e: dataout_d = 16'h0086;
         10'h35f: dataout_d = 16'h0068;
         10'h360: dataout_d = 16'h0085;
         10'h361: dataout_d = 16'h0083;
         10'h362: dataout_d = 16'h0068;
         10'h363: dataout_d = 16'h0085;
         10'h364: dataout_d = 16'h0084;
         10'h365: dataout_d = 16'h00a0;
         10'h366: dataout_d = 16'h0001;
         10'h367: dataout_d = 16'h00b1;
         10'h368: dataout_d = 16'h0083;
         10'h369: dataout_d = 16'h00e6;
         10'h36a: dataout_d = 16'h0083;
         10'h36b: dataout_d = 16'h00d0;
         10'h36c: dataout_d = 16'h0002;
         10'h36d: dataout_d = 16'h00e6;
         10'h36e: dataout_d = 16'h0084;
         10'h36f: dataout_d = 16'h0009;
         10'h370: dataout_d = 16'h0000;
         10'h371: dataout_d = 16'h00f0;
         10'h372: dataout_d = 16'h0006;
         10'h373: dataout_d = 16'h0020;
         10'h374: dataout_d = 16'hff97;
         10'h375: dataout_d = 16'hffff;
         10'h376: dataout_d = 16'h004c;
         10'h377: dataout_d = 16'hff65;
         10'h378: dataout_d = 16'hffff;
         10'h379: dataout_d = 16'h00e6;
         10'h37a: dataout_d = 16'h0083;
         10'h37b: dataout_d = 16'h00d0;
         10'h37c: dataout_d = 16'h0002;
         10'h37d: dataout_d = 16'h00e6;
         10'h37e: dataout_d = 16'h0084;
         10'h37f: dataout_d = 16'h00a4;
         10'h380: dataout_d = 16'h0086;
         10'h381: dataout_d = 16'h006c;
         10'h382: dataout_d = 16'h0083;
         10'h383: dataout_d = 16'h0000;
         10'h384: dataout_d = 16'h0048;
         10'h385: dataout_d = 16'h004a;
         10'h386: dataout_d = 16'h004a;
         10'h387: dataout_d = 16'h004a;
         10'h388: dataout_d = 16'h004a;
         10'h389: dataout_d = 16'h0020;
         10'h38a: dataout_d = 16'hff8d;
         10'h38b: dataout_d = 16'hffff;
         10'h38c: dataout_d = 16'h0068;
         10'h38d: dataout_d = 16'h0029;
         10'h38e: dataout_d = 16'h000f;
         10'h38f: dataout_d = 16'h00c9;
         10'h390: dataout_d = 16'h000a;
         10'h391: dataout_d = 16'h0090;
         10'h392: dataout_d = 16'h0002;
         10'h393: dataout_d = 16'h0069;
         10'h394: dataout_d = 16'h0006;
         10'h395: dataout_d = 16'h0069;
         10'h396: dataout_d = 16'h0030;
         10'h397: dataout_d = 16'h0048;
         10'h398: dataout_d = 16'h00ad;
         10'h399: dataout_d = 16'hfff8;
         10'h39a: dataout_d = 16'hfffa;
         10'h39b: dataout_d = 16'h004a;
         10'h39c: dataout_d = 16'h004a;
         10'h39d: dataout_d = 16'h0090;
         10'h39e: dataout_d = 16'hfff9;
         10'h39f: dataout_d = 16'h0068;
         10'h3a0: dataout_d = 16'h008d;
         10'h3a1: dataout_d = 16'hfff9;
         10'h3a2: dataout_d = 16'hfffa;
         10'h3a3: dataout_d = 16'h0060;
         10'h3a4: dataout_d = 16'h0086;
         10'h3a5: dataout_d = 16'h0085;
         10'h3a6: dataout_d = 16'h00a6;
         10'h3a7: dataout_d = 16'h0081;
         10'h3a8: dataout_d = 16'h0095;
         10'h3a9: dataout_d = 16'h0041;
         10'h3aa: dataout_d = 16'h00e8;
         10'h3ab: dataout_d = 16'h008a;
         10'h3ac: dataout_d = 16'h0029;
         10'h3ad: dataout_d = 16'h003f;
         10'h3ae: dataout_d = 16'h0085;
         10'h3af: dataout_d = 16'h0081;
         10'h3b0: dataout_d = 16'h00a6;
         10'h3b1: dataout_d = 16'h0085;
         10'h3b2: dataout_d = 16'h0060;
         10'h3b3: dataout_d = 16'h0040;
         10'h3b4: dataout_d = 16'h0000;
         10'h3b5: dataout_d = 16'h0000;
         10'h3b6: dataout_d = 16'h0000;
         10'h3b7: dataout_d = 16'h0000;
         10'h3b8: dataout_d = 16'h0000;
         10'h3b9: dataout_d = 16'h0000;
         10'h3ba: dataout_d = 16'h0000;
         10'h3bb: dataout_d = 16'h0000;
         10'h3bc: dataout_d = 16'h0000;
         10'h3bd: dataout_d = 16'h0000;
         10'h3be: dataout_d = 16'h0000;
         10'h3bf: dataout_d = 16'h0000;
         10'h3c0: dataout_d = 16'h0000;
         10'h3c1: dataout_d = 16'h0000;
         10'h3c2: dataout_d = 16'h0000;
         10'h3c3: dataout_d = 16'h0000;
         10'h3c4: dataout_d = 16'h0000;
         10'h3c5: dataout_d = 16'h0000;
         10'h3c6: dataout_d = 16'h0000;
         10'h3c7: dataout_d = 16'h0000;
         10'h3c8: dataout_d = 16'h0000;
         10'h3c9: dataout_d = 16'h0000;
         10'h3ca: dataout_d = 16'h0000;
         10'h3cb: dataout_d = 16'h0000;
         10'h3cc: dataout_d = 16'h0000;
         10'h3cd: dataout_d = 16'h0000;
         10'h3ce: dataout_d = 16'h0000;
         10'h3cf: dataout_d = 16'h0000;
         10'h3d0: dataout_d = 16'h0000;
         10'h3d1: dataout_d = 16'h0000;
         10'h3d2: dataout_d = 16'h0000;
         10'h3d3: dataout_d = 16'h0000;
         10'h3d4: dataout_d = 16'h0000;
         10'h3d5: dataout_d = 16'h0000;
         10'h3d6: dataout_d = 16'h0000;
         10'h3d7: dataout_d = 16'h0000;
         10'h3d8: dataout_d = 16'h0000;
         10'h3d9: dataout_d = 16'h0000;
         10'h3da: dataout_d = 16'h0000;
         10'h3db: dataout_d = 16'h0000;
         10'h3dc: dataout_d = 16'h0000;
         10'h3dd: dataout_d = 16'h0000;
         10'h3de: dataout_d = 16'h0000;
         10'h3df: dataout_d = 16'h0000;
         10'h3e0: dataout_d = 16'h004c;
         10'h3e1: dataout_d = 16'hff35;
         10'h3e2: dataout_d = 16'hffff;
         10'h3e3: dataout_d = 16'h0000;
         10'h3e4: dataout_d = 16'h0000;
         10'h3e5: dataout_d = 16'h0000;
         10'h3e6: dataout_d = 16'h0000;
         10'h3e7: dataout_d = 16'h0000;
         10'h3e8: dataout_d = 16'h0000;
         10'h3e9: dataout_d = 16'h0000;
         10'h3ea: dataout_d = 16'h0000;
         10'h3eb: dataout_d = 16'h0000;
         10'h3ec: dataout_d = 16'h0000;
         10'h3ed: dataout_d = 16'h0000;
         10'h3ee: dataout_d = 16'h004c;
         10'h3ef: dataout_d = 16'hff97;
         10'h3f0: dataout_d = 16'hffff;
         10'h3f1: dataout_d = 16'h0000;
         10'h3f2: dataout_d = 16'h0000;
         10'h3f3: dataout_d = 16'h0000;
         10'h3f4: dataout_d = 16'h0000;
         10'h3f5: dataout_d = 16'h0000;
         10'h3f6: dataout_d = 16'h0000;
         10'h3f7: dataout_d = 16'h0000;
         10'h3f8: dataout_d = 16'h0000;
         10'h3f9: dataout_d = 16'h0000;
         10'h3fa: dataout_d = 16'hffb3;
         10'h3fb: dataout_d = 16'hffff;
         10'h3fc: dataout_d = 16'hfd80;
         10'h3fd: dataout_d = 16'hffff;
         10'h3fe: dataout_d = 16'hffb3;
         10'h3ff: dataout_d = 16'hffff;

	 default:
	   begin
	     dataout_d = 16'hxxxx;
	   end
       endcase
     end

endmodule
